library IEEE; use IEEE.STD_LOGIC_1164.all; use IEEE.NUMERIC_STD.all;

entity main is
port(
	clk, data_in, rst_n : in STD_LOGIC;
	stored_val : out STD_LOGIC_VECTOR(7 downto 0);
	counter_out : out UNSIGNED(3 downto 0)

);
end entity main; 

architecture synth of main is
--signal declaration
CONSTANT clk_freq : integer := 25_000_000; --ENTER FREQUENCY HERE!
CONSTANT baud_rate : integer := 9600; --ENTER BAUDRATE HERE!
CONSTANT bit_time : integer := clk_freq/baud_rate;
signal reg : STD_LOGIC_VECTOR(7 downto 0) := (others=>'0');
signal counter : UNSIGNED(3 downto 0);
signal timer : UNSIGNED(11 downto 0);
type statetype is (IDLEREAD, IDLEWAIT, OPREAD, OPWAIT, STOPWAIT);
signal state : statetype;
begin
--main control process
process(clk)
begin
if(rising_edge(clk)) then
	--reset conditions
	if(rst_n = '0') then
		state <= IDLEREAD;
		counter <= (others => '0');
	else
	--initialization
	if(state = IDLEREAD and data_in = '0') then
		state <= IDLEWAIT;
		counter <= (others => '0');
	elsif(state = IDLEWAIT) then
	--initial waiting (1.5 times)
	if(timer = bit_time + bit_time/2) then
		state <= OPREAD;
	end if; --end initial waiting
	end if; --end initialization if
	--reading normal data
	if(state = OPREAD) then
		state <= OPWAIT;
		counter <= counter + 1;
	end if;
	--waiting between normal data inputs
	if(state = OPWAIT) then
		if(timer = bit_time and counter /= 8) then		
		state <= OPREAD;
		--ending condition, triggers after the last bit has been inputted
		elsif(counter = 8 and state = OPWAIT) then
			state <= STOPWAIT;
		end if;
	end if;
	--stop condition
	if(state = STOPWAIT) then
		if(timer = bit_time) then
			state <= IDLEREAD;
		end if;
	end if;
	
	end if;
end if;
end process;

--timer process
process(clk) 
begin
if(rising_edge(clk)) then
if(rst_n='1') then
	if(state = IDLEWAIT or state = OPWAIT or state = STOPWAIT) then
		timer <= timer + 1;
	else
		timer <= (others => '0');
	end if;
else
	timer <= (others => '0');
end if;
end if;
end process;

--reader process
process(clk)
begin
if(rising_edge(clk)) then
	if(state = OPREAD) then
		reg <= data_in & reg(7 downto 1);

	end if;
	if(state = IDLEREAD) then
		reg <= (others=>'0');
	end if;
end if;
end process;

--outputs
stored_val <= reg;
counter_out <= counter;
end architecture synth;